LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY LED_16 IS
	PORT(A:INTEGER RANGE 0 TO 15;
		LED7:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END LED_16;
ARCHITECTURE ONE OF LED_16 IS
BEGIN
	PROCESS(A)
	BEGIN
	CASE A IS
		WHEN 0 => LED7 <= "00111111";
		WHEN 1 => LED7 <= "00000110";
		WHEN 2 => LED7 <= "01011011";
		WHEN 3 => LED7 <= "01001111";
		WHEN 4 => LED7 <= "01100110";
		WHEN 5 => LED7 <= "01101101";
		WHEN 6 => LED7 <= "01111101";
		WHEN 7 => LED7 <= "00000111";
		WHEN 8 => LED7 <= "01111111";
		WHEN 9 => LED7 <= "01101111";
		WHEN 10 => LED7 <= "01110111";
		WHEN 11 => LED7 <= "01111100";
		WHEN 12 => LED7 <= "00111001";
		WHEN 13 => LED7 <= "01011110";
		WHEN 14 => LED7 <= "01111001";
		WHEN 15 => LED7 <= "01110001";
		WHEN OTHERS => NULL;
	END CASE;
END PROCESS;
END ONE;
	