LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY COUNTER_TOP IS
	PORT(CLK,EN0:IN STD_LOGIC;
		COUT4:OUT STD_LOGIC;
		HEX0,HEX1:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));

END COUNTER_TOP;
ARCHITECTURE ONE OF COUNTER_TOP IS

COMPONENT Counter_lsl 
PORT(CLK,EN:IN STD_LOGIC;
		COUT:OUT STD_LOGIC;
		Q:BUFFER INTEGER RANGE 0 TO 15);
END COMPONENT;

COMPONENT LED_16
PORT(A:INTEGER RANGE 0 TO 15;
		LED7:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT Timer_lsl
port(CLKIN	:in std_logic;   
	 CLKOUT	:out std_logic
);
END COMPONENT;

SIGNAL CLK1,COUT0:STD_LOGIC;
SIGNAL Q0,Q1:INTEGER RANGE 0 TO 15;

BEGIN
U1:Timer_lsl PORT MAP (CLKIN => CLK,CLKOUT => CLK1);
U2:Counter_lsl PORT MAP (CLK => CLK1,EN => EN0, COUT => COUT0,Q=>Q0);
U3:Counter_lsl PORT MAP (CLK => CLK1,EN =>COUT0, COUT => COUT4,Q=>Q1);
U4:LED_16 PORT MAP(A => Q0,LED7 => HEX0);
U5:LED_16 PORT MAP(A => Q1,LED7 => HEX1);
END ONE;